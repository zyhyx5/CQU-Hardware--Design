`include "../my_mips.svh"
`include "../define.svh"

module exception (
    input  logic            rst,
    input  exception_sign_t exception_sign,
    output exception_data_t exception_data

);




endmodule
